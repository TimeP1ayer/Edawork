//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sun Dec 24 20:43:40 2023
// Version: v11.9 SP1 11.9.1.0
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// ex4511_161
module ex4511_161(
    // Inputs
    CP,
    Dn,
    LE,
    // Outputs
    Seg,
    TC
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        CP;
input  [3:0] Dn;
input        LE;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0] Seg;
output       TC;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         CP;
wire   [3:0] Dn;
wire   [3:0] HC161_0_Qn;
wire   [1:1] HC161_0_Qn1to1;
wire   [3:3] HC161_0_Qn3to3;
wire         LE;
wire         NAND2_0_Y;
wire   [7:0] Seg_net_0;
wire         TC_net_0;
wire   [7:0] Seg_net_1;
wire         TC_net_1;
wire   [0:0] Qn_slice_0;
wire   [2:2] Qn_slice_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         VCC_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net = 1'b1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Seg_net_1 = Seg_net_0;
assign Seg[7:0]  = Seg_net_1;
assign TC_net_1  = TC_net_0;
assign TC        = TC_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign HC161_0_Qn1to1[1] = HC161_0_Qn[1:1];
assign HC161_0_Qn3to3[3] = HC161_0_Qn[3:3];
assign Qn_slice_0[0]     = HC161_0_Qn[0:0];
assign Qn_slice_1[2]     = HC161_0_Qn[2:2];
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------HC161
HC161 HC161_0(
        // Inputs
        .CP  ( CP ),
        .CEP ( VCC_net ),
        .CET ( VCC_net ),
        .MRN ( NAND2_0_Y ),
        .PEN ( VCC_net ),
        .Dn  ( Dn ),
        // Outputs
        .Qn  ( HC161_0_Qn ),
        .TC  ( TC_net_0 ) 
        );

//--------hc4511
hc4511 hc4511_0(
        // Inputs
        .LE   ( LE ),
        .BI_N ( VCC_net ),
        .LT_N ( VCC_net ),
        .A    ( HC161_0_Qn ),
        // Outputs
        .Seg  ( Seg_net_0 ) 
        );

//--------NAND2
NAND2 NAND2_0(
        // Inputs
        .A ( HC161_0_Qn3to3 ),
        .B ( HC161_0_Qn1to1 ),
        // Outputs
        .Y ( NAND2_0_Y ) 
        );


endmodule
