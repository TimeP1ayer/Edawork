//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Wed Jan 03 14:04:45 2024
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// ex161ex4511
module ex161ex4511(
    // Inputs
    CP,
    Dn,
    MRN,
    // Outputs
    Seg
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        CP;
input  [3:0] Dn;
input        MRN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0] Seg;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         CP;
wire   [3:0] Dn;
wire         MRN;
wire   [3:0] Qn;
wire   [7:0] Seg_net_0;
wire   [7:0] Seg_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         VCC_net;
wire         GND_net;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net = 1'b1;
assign GND_net = 1'b0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Seg_net_1 = Seg_net_0;
assign Seg[7:0]  = Seg_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------HC161
HC161 HC161_0(
        // Inputs
        .CP  ( CP ),
        .CEP ( VCC_net ),
        .CET ( VCC_net ),
        .MRN ( MRN ),
        .PEN ( VCC_net ),
        .Dn  ( Dn ),
        // Outputs
        .Qn  ( Qn ),
        .TC  (  ) 
        );

//--------hc4511
hc4511 hc4511_0(
        // Inputs
        .LE   ( GND_net ),
        .BI_N ( VCC_net ),
        .LT_N ( VCC_net ),
        .A    ( Qn ),
        // Outputs
        .Seg  ( Seg_net_0 ) 
        );


endmodule
