///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: hc2831.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::ProASIC3> <Die::A3P060> <Package::100 VQFP>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module hc2831( port1, port2, port3, port4 );
input port1, port2;
output port3;
inout port4;

//<statements>

endmodule

